//=======================================================
// ECE3400 Fall 2017
// Lab 3: Template ROM module
//
// Top-level skeleton from Terasic
// Modified by Claire Chen for ECE3400 Fall 2017
//=======================================================

module G5_783_ROM(	
	input [8:0] addr,
	input clk,
	output reg [7:0] q
);

    //=======================================================
    //  REG/WIRE declarations
    //=======================================================
	 reg [7:0] sin[159:0];
	 
	 initial begin
		sin[0]  <= 8'b10000000;
		sin[1]  <= 8'b10000101;
		sin[2]  <= 8'b10001010;
		sin[3]  <= 8'b10001111;
		sin[4]  <= 8'b10010100;
		sin[5]  <= 8'b10011000;
		sin[6]  <= 8'b10011101;
		sin[7]  <= 8'b10100010;
		sin[8]  <= 8'b10100111;
		sin[9]  <= 8'b10101100;
		sin[10] <= 8'b10110000;
		sin[11] <= 8'b10110101;
		sin[12] <= 8'b10111010;
		sin[13] <= 8'b10111110;
		sin[14] <= 8'b11000010;
		sin[15] <= 8'b11000111;
		sin[16] <= 8'b11001011;
		sin[17] <= 8'b11001111;
		sin[18] <= 8'b11010011;
		sin[19] <= 8'b11010110;
		sin[20] <= 8'b11011010;
		sin[21] <= 8'b11011101;
		sin[22] <= 8'b11100001;
		sin[23] <= 8'b11100100;
		sin[24] <= 8'b11100111;
		sin[25] <= 8'b11101010;
		sin[26] <= 8'b11101100;
		sin[27] <= 8'b11101111;
		sin[28] <= 8'b11110001;
		sin[29] <= 8'b11110100;
		sin[30] <= 8'b11110101;
		sin[31] <= 8'b11110111;
		sin[32] <= 8'b11111001;
		sin[33] <= 8'b11111010;
		sin[34] <= 8'b11111100;
		sin[35] <= 8'b11111101;
		sin[36] <= 8'b11111110;
		sin[37] <= 8'b11111110;
		sin[38] <= 8'b11111111;
		sin[39] <= 8'b11111111;
		sin[40] <= 8'b11111111;
		sin[41] <= 8'b11111111;
		sin[42] <= 8'b11111111;
		sin[43] <= 8'b11111110;
		sin[44] <= 8'b11111101;
		sin[45] <= 8'b11111100;
		sin[46] <= 8'b11111011;
		sin[47] <= 8'b11111010;
		sin[48] <= 8'b11111000;
		sin[49] <= 8'b11110111;
		sin[50] <= 8'b11110101;
		sin[51] <= 8'b11110011;
		sin[52] <= 8'b11110001;
		sin[53] <= 8'b11101110;
		sin[54] <= 8'b11101100;
		sin[55] <= 8'b11101001;
		sin[56] <= 8'b11100110;
		sin[57] <= 8'b11100011;
		sin[58] <= 8'b11100000;
		sin[59] <= 8'b11011100;
		sin[60] <= 8'b11011001;
		sin[61] <= 8'b11010101;
		sin[62] <= 8'b11010001;
		sin[63] <= 8'b11001110;
		sin[64] <= 8'b11001010;
		sin[65] <= 8'b11000101;
		sin[66] <= 8'b11000001;
		sin[67] <= 8'b10111101;
		sin[68] <= 8'b10111000;
		sin[69] <= 8'b10110100;
		sin[70] <= 8'b10101111;
		sin[71] <= 8'b10101010;
		sin[72] <= 8'b10100110;
		sin[73] <= 8'b10100001;
		sin[74] <= 8'b10011100;
		sin[75] <= 8'b10010111;
		sin[76] <= 8'b10010010;
		sin[77] <= 8'b10001101;
		sin[78] <= 8'b10001000;
		sin[79] <= 8'b10000011;
		sin[80] <= 8'b01111110;
		sin[81] <= 8'b01111001;
		sin[82] <= 8'b01110100;
		sin[83] <= 8'b01101111;
		sin[84] <= 8'b01101010;
		sin[85] <= 8'b01100101;
		sin[86] <= 8'b01100000;
		sin[87] <= 8'b01011011;
		sin[88] <= 8'b01010111;
		sin[89] <= 8'b01010010;
		sin[90] <= 8'b01001101;
		sin[91] <= 8'b01001001;
		sin[92] <= 8'b01000100;
		sin[93] <= 8'b01000000;
		sin[94] <= 8'b00111011;
		sin[95] <= 8'b00110111;
		sin[96] <= 8'b00110011;
		sin[97] <= 8'b00101111;
		sin[98] <= 8'b00101011;
		sin[99] <= 8'b00101000;
		sin[100] <= 8'b00100100;
		sin[101] <= 8'b00100001;
		sin[102] <= 8'b00011101;
		sin[103] <= 8'b00011010;
		sin[104] <= 8'b00010111;
		sin[105] <= 8'b00010100;
		sin[106] <= 8'b00010010;
		sin[107] <= 8'b00001111;
		sin[108] <= 8'b00001101;
		sin[109] <= 8'b00001011;
		sin[110] <= 8'b00001001;
		sin[111] <= 8'b00000111;
		sin[112] <= 8'b00000110;
		sin[113] <= 8'b00000100;
		sin[114] <= 8'b00000011;
		sin[115] <= 8'b00000010;
		sin[116] <= 8'b00000001;
		sin[117] <= 8'b00000001;
		sin[118] <= 8'b00000000;
		sin[119] <= 8'b00000000;
		sin[120] <= 8'b00000000;
		sin[121] <= 8'b00000000;
		sin[122] <= 8'b00000001;
		sin[123] <= 8'b00000001;
		sin[124] <= 8'b00000010;
		sin[125] <= 8'b00000011;
		sin[126] <= 8'b00000100;
		sin[127] <= 8'b00000101;
		sin[128] <= 8'b00000111;
		sin[129] <= 8'b00001001;
		sin[130] <= 8'b00001011;
		sin[131] <= 8'b00001101;
		sin[132] <= 8'b00001111;
		sin[133] <= 8'b00010001;
		sin[134] <= 8'b00010100;
		sin[135] <= 8'b00010111;
		sin[136] <= 8'b00011010;
		sin[137] <= 8'b00011101;
		sin[138] <= 8'b00100000;
		sin[139] <= 8'b00100100;
		sin[140] <= 8'b00100111;
		sin[141] <= 8'b00101011;
		sin[142] <= 8'b00101111;
		sin[143] <= 8'b00110011;
		sin[144] <= 8'b00110111;
		sin[145] <= 8'b00111011;
		sin[146] <= 8'b00111111;
		sin[147] <= 8'b01000011;
		sin[148] <= 8'b01001000;
		sin[149] <= 8'b01001101;
		sin[150] <= 8'b01010001;
		sin[151] <= 8'b01010110;
		sin[152] <= 8'b01011011;
		sin[153] <= 8'b01011111;
		sin[154] <= 8'b01100100;
		sin[155] <= 8'b01101001;
		sin[156] <= 8'b01101110;
		sin[157] <= 8'b01110011;
		sin[158] <= 8'b01111000;
		sin[159] <= 8'b01111101;
	 end
	 
    //=======================================================
    //  Structural coding
    //=======================================================
	 always @(posedge clk) begin
		q <= sin[addr];
	 end
	 
endmodule