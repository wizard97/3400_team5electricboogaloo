//=======================================================
// ECE3400 Fall 2017
// Lab 3: Template top-level module
//
// Top-level skeleton from Terasic
// Modified by Claire Chen for ECE3400 Fall 2017
//=======================================================

`define ONE_SEC 25000000

module DE0_NANO(

	//////////// CLOCK //////////
	CLOCK_50,

	//////////// LED //////////
	//LED,

	//////////// KEY //////////
	KEY,

	//////////// SW //////////
	//SW,

	//////////// GPIO_0, GPIO_0 connect to GPIO Default //////////
	GPIO_0_D,
	//GPIO_0_IN,

	//////////// GPIO_0, GPIO_1 connect to GPIO Default //////////
	//GPIO_1_D,
	//GPIO_1_IN,
	
//	GPIO_2_IN,
//	GPIO_3_IN,
//	GPIO_4_IN,
//	GPIO_5_IN,
//	GPIO_6_IN,
//	GPIO_7_IN,
//	GPIO_8_IN,
//	GPIO_9_IN
);

	  //=======================================================
	 //  PARAMETER declarations
	 //=======================================================

	 localparam COUNT = 25000000/440/2; // one second in 25MHz clock cycles
	 
	 //=======================================================
	 //  PORT declarations
	 //=======================================================

	 //////////// CLOCK //////////
	 input 		          		CLOCK_50;

	 //////////// LED //////////
	 //output		     [7:0]		LED;

	 /////////// KEY //////////
	 input 		     [1:0]		KEY;

	 //////////// SW //////////
	 //input 		     [3:0]		SW;

	 //////////// GPIO_0, GPIO_0 connect to GPIO Default //////////
	 inout 		    [33:0]		GPIO_0_D;
	 //input 		     [1:0]		GPIO_0_IN;

	 //////////// GPIO_0, GPIO_1 connect to GPIO Default //////////
	 //inout 		    [33:0]		GPIO_1_D;
	 //input 		     [1:0]		GPIO_1_IN;
	 
//	 input			  [1:0]		GPIO_2_IN;
//	 input			  [1:0]		GPIO_3_IN;
//	 input			  [1:0]		GPIO_4_IN;
//	 input			  [1:0]		GPIO_5_IN;
//	 input			  [1:0]		GPIO_6_IN;
//	 input			  [1:0]		GPIO_7_IN;
//	 input			  [1:0]		GPIO_8_IN;
//	 input			  [1:0]		GPIO_9_IN;

    //=======================================================

    //=======================================================
    //  REG/WIRE declarations
    //=======================================================
    reg         CLOCK_25;
    wire        reset; // active high reset signal 

//    wire [9:0]  PIXEL_COORD_X; // current x-coord from VGA driver
//    wire [9:0]  PIXEL_COORD_Y; // current y-coord from VGA driver
//    wire [7:0]  PIXEL_COLOR;   // input 8-bit pixel color for current coords
//	 
//	 reg [24:0] led_counter; // timer to keep track of when to toggle LED
//	 reg 			led_state;   // 1 is on, 0 is off

		reg  [6:0] counter;
		reg  [9:0] addr;
		wire [7:0] q;
//	 
    // Module outputs coordinates of next pixel to be written onto screen
//    VGA_DRIVER driver(
//		  .RESET(reset),
//        .CLOCK(CLOCK_25),
//        .PIXEL_COLOR_IN(PIXEL_COLOR),
//        .PIXEL_X(PIXEL_COORD_X),
//        .PIXEL_Y(PIXEL_COORD_Y),
//        .PIXEL_COLOR_OUT({GPIO_0_D[9],GPIO_0_D[11],GPIO_0_D[13],GPIO_0_D[15],GPIO_0_D[17],GPIO_0_D[19],GPIO_0_D[21],GPIO_0_D[23]}),
//        .H_SYNC_NEG(GPIO_0_D[7]),
//        .V_SYNC_NEG(GPIO_0_D[5])
//    );
//	 

		SINE_ROM sine_table(
			.addr(addr),
			.clk(CLOCK_25),
			.q(q)
		);
		
		assign GPIO_0_D[0] = q[0];
		assign GPIO_0_D[1] = q[1];
		assign GPIO_0_D[2] = q[2];
		assign GPIO_0_D[3] = q[3];
		assign GPIO_0_D[4] = q[4];
		assign GPIO_0_D[5] = q[5];
		assign GPIO_0_D[6] = q[6];
		assign GPIO_0_D[7] = q[7];
		
	 assign reset = ~KEY[0]; // reset when KEY0 is pressed
//	 
//	 assign PIXEL_COLOR = 8'b000_111_00; // Green
//	 assign LED[0] = led_state;
	 
    //=======================================================
    //  Structural coding
    //=======================================================
 
	 // Generate 25MHz clock for VGA, FPGA has 50 MHz clock
    always @ (posedge CLOCK_50) begin
        CLOCK_25 <= ~CLOCK_25; 
    end // always @ (posedge CLOCK_50)
	
	 // Simple state machine to toggle square wave every one second
	 always @ (posedge CLOCK_25) begin
		  if (reset) begin
				counter   <= 90;
				addr      <= 0;
		  end
		  
		  else if (counter == 0) begin
				counter   <= 90;
				if (addr == 632) begin
					addr <= 0;
				end
				else begin
					addr      <= addr + 1;
				end
		  end
		  /*if (led_counter == ONE_SEC) begin
				led_state   <= ~led_state;
				led_counter <= 25'b0;
		  end*/
		  else begin	
				//led_state   <= led_state;
				counter	 <= counter - 1;
		  end // always @ (posedge CLOCK_25)
		  
		  //sin <= q;
	 end
	 

endmodule
