//=======================================================
// ECE3400 Fall 2017
// Lab 3: Template ROM module
//
// Top-level skeleton from Terasic
// Modified by Claire Chen for ECE3400 Fall 2017
//=======================================================

module G4_392_ROM(	
	input [9:0] addr,
	input clk,
	output reg [7:0] q
);

    //=======================================================
    //  REG/WIRE declarations
    //=======================================================
	 reg [7:0] sin[318:0];
	 
	 initial begin
		sin[0]  <= 8'b10000000;
		sin[1]  <= 8'b10000010;
		sin[2]  <= 8'b10000101;
		sin[3]  <= 8'b10000111;
		sin[4]  <= 8'b10001010;
		sin[5]  <= 8'b10001100;
		sin[6]  <= 8'b10001111;
		sin[7]  <= 8'b10010001;
		sin[8]  <= 8'b10010100;
		sin[9]  <= 8'b10010110;
		sin[10] <= 8'b10011000;
		sin[11] <= 8'b10011011;
		sin[12] <= 8'b10011101;
		sin[13] <= 8'b10100000;
		sin[14] <= 8'b10100010;
		sin[15] <= 8'b10100101;
		sin[16] <= 8'b10100111;
		sin[17] <= 8'b10101001;
		sin[18] <= 8'b10101100;
		sin[19] <= 8'b10101110;
		sin[20] <= 8'b10110000;
		sin[21] <= 8'b10110011;
		sin[22] <= 8'b10110101;
		sin[23] <= 8'b10110111;
		sin[24] <= 8'b10111010;
		sin[25] <= 8'b10111100;
		sin[26] <= 8'b10111110;
		sin[27] <= 8'b11000000;
		sin[28] <= 8'b11000010;
		sin[29] <= 8'b11000100;
		sin[30] <= 8'b11000111;
		sin[31] <= 8'b11001001;
		sin[32] <= 8'b11001011;
		sin[33] <= 8'b11001101;
		sin[34] <= 8'b11001111;
		sin[35] <= 8'b11010001;
		sin[36] <= 8'b11010011;
		sin[37] <= 8'b11010100;
		sin[38] <= 8'b11010110;
		sin[39] <= 8'b11011000;
		sin[40] <= 8'b11011010;
		sin[41] <= 8'b11011100;
		sin[42] <= 8'b11011101;
		sin[43] <= 8'b11011111;
		sin[44] <= 8'b11100001;
		sin[45] <= 8'b11100010;
		sin[46] <= 8'b11100100;
		sin[47] <= 8'b11100101;
		sin[48] <= 8'b11100111;
		sin[49] <= 8'b11101000;
		sin[50] <= 8'b11101010;
		sin[51] <= 8'b11101011;
		sin[52] <= 8'b11101100;
		sin[53] <= 8'b11101110;
		sin[54] <= 8'b11101111;
		sin[55] <= 8'b11110000;
		sin[56] <= 8'b11110001;
		sin[57] <= 8'b11110010;
		sin[58] <= 8'b11110100;
		sin[59] <= 8'b11110101;
		sin[60] <= 8'b11110101;
		sin[61] <= 8'b11110110;
		sin[62] <= 8'b11110111;
		sin[63] <= 8'b11111000;
		sin[64] <= 8'b11111001;
		sin[65] <= 8'b11111010;
		sin[66] <= 8'b11111010;
		sin[67] <= 8'b11111011;
		sin[68] <= 8'b11111100;
		sin[69] <= 8'b11111100;
		sin[70] <= 8'b11111101;
		sin[71] <= 8'b11111101;
		sin[72] <= 8'b11111110;
		sin[73] <= 8'b11111110;
		sin[74] <= 8'b11111110;
		sin[75] <= 8'b11111110;
		sin[76] <= 8'b11111111;
		sin[77] <= 8'b11111111;
		sin[78] <= 8'b11111111;
		sin[79] <= 8'b11111111;
		sin[80] <= 8'b11111111;
		sin[81] <= 8'b11111111;
		sin[82] <= 8'b11111111;
		sin[83] <= 8'b11111111;
		sin[84] <= 8'b11111111;
		sin[85] <= 8'b11111110;
		sin[86] <= 8'b11111110;
		sin[87] <= 8'b11111110;
		sin[88] <= 8'b11111101;
		sin[89] <= 8'b11111101;
		sin[90] <= 8'b11111100;
		sin[91] <= 8'b11111100;
		sin[92] <= 8'b11111011;
		sin[93] <= 8'b11111011;
		sin[94] <= 8'b11111010;
		sin[95] <= 8'b11111001;
		sin[96] <= 8'b11111000;
		sin[97] <= 8'b11111000;
		sin[98] <= 8'b11110111;
		sin[99] <= 8'b11110110;
		sin[100] <= 8'b11110101;
		sin[101] <= 8'b11110100;
		sin[102] <= 8'b11110011;
		sin[103] <= 8'b11110010;
		sin[104] <= 8'b11110001;
		sin[105] <= 8'b11110000;
		sin[106] <= 8'b11101110;
		sin[107] <= 8'b11101101;
		sin[108] <= 8'b11101100;
		sin[109] <= 8'b11101010;
		sin[110] <= 8'b11101001;
		sin[111] <= 8'b11101000;
		sin[112] <= 8'b11100110;
		sin[113] <= 8'b11100101;
		sin[114] <= 8'b11100011;
		sin[115] <= 8'b11100001;
		sin[116] <= 8'b11100000;
		sin[117] <= 8'b11011110;
		sin[118] <= 8'b11011100;
		sin[119] <= 8'b11011011;
		sin[120] <= 8'b11011001;
		sin[121] <= 8'b11010111;
		sin[122] <= 8'b11010101;
		sin[123] <= 8'b11010011;
		sin[124] <= 8'b11010001;
		sin[125] <= 8'b11010000;
		sin[126] <= 8'b11001110;
		sin[127] <= 8'b11001100;
		sin[128] <= 8'b11001010;
		sin[129] <= 8'b11000111;
		sin[130] <= 8'b11000101;
		sin[131] <= 8'b11000011;
		sin[132] <= 8'b11000001;
		sin[133] <= 8'b10111111;
		sin[134] <= 8'b10111101;
		sin[135] <= 8'b10111011;
		sin[136] <= 8'b10111000;
		sin[137] <= 8'b10110110;
		sin[138] <= 8'b10110100;
		sin[139] <= 8'b10110001;
		sin[140] <= 8'b10101111;
		sin[141] <= 8'b10101101;
		sin[142] <= 8'b10101010;
		sin[143] <= 8'b10101000;
		sin[144] <= 8'b10100110;
		sin[145] <= 8'b10100011;
		sin[146] <= 8'b10100001;
		sin[147] <= 8'b10011110;
		sin[148] <= 8'b10011100;
		sin[149] <= 8'b10011010;
		sin[150] <= 8'b10010111;
		sin[151] <= 8'b10010101;
		sin[152] <= 8'b10010010;
		sin[153] <= 8'b10010000;
		sin[154] <= 8'b10001101;
		sin[155] <= 8'b10001011;
		sin[156] <= 8'b10001000;
		sin[157] <= 8'b10000110;
		sin[158] <= 8'b10000011;
		sin[159] <= 8'b10000001;
		sin[160] <= 8'b01111110;
		sin[161] <= 8'b01111100;
		sin[162] <= 8'b01111001;
		sin[163] <= 8'b01110111;
		sin[164] <= 8'b01110100;
		sin[165] <= 8'b01110010;
		sin[166] <= 8'b01101111;
		sin[167] <= 8'b01101101;
		sin[168] <= 8'b01101010;
		sin[169] <= 8'b01101000;
		sin[170] <= 8'b01100101;
		sin[171] <= 8'b01100011;
		sin[172] <= 8'b01100000;
		sin[173] <= 8'b01011110;
		sin[174] <= 8'b01011011;
		sin[175] <= 8'b01011001;
		sin[176] <= 8'b01010111;
		sin[177] <= 8'b01010100;
		sin[178] <= 8'b01010010;
		sin[179] <= 8'b01010000;
		sin[180] <= 8'b01001101;
		sin[181] <= 8'b01001011;
		sin[182] <= 8'b01001001;
		sin[183] <= 8'b01000110;
		sin[184] <= 8'b01000100;
		sin[185] <= 8'b01000010;
		sin[186] <= 8'b01000000;
		sin[187] <= 8'b00111110;
		sin[188] <= 8'b00111011;
		sin[189] <= 8'b00111001;
		sin[190] <= 8'b00110111;
		sin[191] <= 8'b00110101;
		sin[192] <= 8'b00110011;
		sin[193] <= 8'b00110001;
		sin[194] <= 8'b00101111;
		sin[195] <= 8'b00101101;
		sin[196] <= 8'b00101011;
		sin[197] <= 8'b00101010;
		sin[198] <= 8'b00101000;
		sin[199] <= 8'b00100110;
		sin[200] <= 8'b00100100;
		sin[201] <= 8'b00100010;
		sin[202] <= 8'b00100001;
		sin[203] <= 8'b00011111;
		sin[204] <= 8'b00011101;
		sin[205] <= 8'b00011100;
		sin[206] <= 8'b00011010;
		sin[207] <= 8'b00011001;
		sin[208] <= 8'b00010111;
		sin[209] <= 8'b00010110;
		sin[210] <= 8'b00010100;
		sin[211] <= 8'b00010011;
		sin[212] <= 8'b00010010;
		sin[213] <= 8'b00010001;
		sin[214] <= 8'b00001111;
		sin[215] <= 8'b00001110;
		sin[216] <= 8'b00001101;
		sin[217] <= 8'b00001100;
		sin[218] <= 8'b00001011;
		sin[219] <= 8'b00001010;
		sin[220] <= 8'b00001001;
		sin[221] <= 8'b00001000;
		sin[222] <= 8'b00000111;
		sin[223] <= 8'b00000110;
		sin[224] <= 8'b00000110;
		sin[225] <= 8'b00000101;
		sin[226] <= 8'b00000100;
		sin[227] <= 8'b00000100;
		sin[228] <= 8'b00000011;
		sin[229] <= 8'b00000011;
		sin[230] <= 8'b00000010;
		sin[231] <= 8'b00000010;
		sin[232] <= 8'b00000001;
		sin[233] <= 8'b00000001;
		sin[234] <= 8'b00000001;
		sin[235] <= 8'b00000000;
		sin[236] <= 8'b00000000;
		sin[237] <= 8'b00000000;
		sin[238] <= 8'b00000000;
		sin[239] <= 8'b00000000;
		sin[240] <= 8'b00000000;
		sin[241] <= 8'b00000000;
		sin[242] <= 8'b00000000;
		sin[243] <= 8'b00000000;
		sin[244] <= 8'b00000001;
		sin[245] <= 8'b00000001;
		sin[246] <= 8'b00000001;
		sin[247] <= 8'b00000010;
		sin[248] <= 8'b00000010;
		sin[249] <= 8'b00000010;
		sin[250] <= 8'b00000011;
		sin[251] <= 8'b00000011;
		sin[252] <= 8'b00000100;
		sin[253] <= 8'b00000101;
		sin[254] <= 8'b00000101;
		sin[255] <= 8'b00000110;
		sin[256] <= 8'b00000111;
		sin[257] <= 8'b00001000;
		sin[258] <= 8'b00001001;
		sin[259] <= 8'b00001010;
		sin[260] <= 8'b00001011;
		sin[261] <= 8'b00001100;
		sin[262] <= 8'b00001101;
		sin[263] <= 8'b00001110;
		sin[264] <= 8'b00001111;
		sin[265] <= 8'b00010000;
		sin[266] <= 8'b00010001;
		sin[267] <= 8'b00010011;
		sin[268] <= 8'b00010100;
		sin[269] <= 8'b00010101;
		sin[270] <= 8'b00010111;
		sin[271] <= 8'b00011000;
		sin[272] <= 8'b00011010;
		sin[273] <= 8'b00011011;
		sin[274] <= 8'b00011101;
		sin[275] <= 8'b00011110;
		sin[276] <= 8'b00100000;
		sin[277] <= 8'b00100010;
		sin[278] <= 8'b00100100;
		sin[279] <= 8'b00100101;
		sin[280] <= 8'b00100111;
		sin[281] <= 8'b00101001;
		sin[282] <= 8'b00101011;
		sin[283] <= 8'b00101101;
		sin[284] <= 8'b00101111;
		sin[285] <= 8'b00110001;
		sin[286] <= 8'b00110011;
		sin[287] <= 8'b00110101;
		sin[288] <= 8'b00110111;
		sin[289] <= 8'b00111001;
		sin[290] <= 8'b00111011;
		sin[291] <= 8'b00111101;
		sin[292] <= 8'b00111111;
		sin[293] <= 8'b01000001;
		sin[294] <= 8'b01000011;
		sin[295] <= 8'b01000110;
		sin[296] <= 8'b01001000;
		sin[297] <= 8'b01001010;
		sin[298] <= 8'b01001101;
		sin[299] <= 8'b01001111;
		sin[300] <= 8'b01010001;
		sin[301] <= 8'b01010100;
		sin[302] <= 8'b01010110;
		sin[303] <= 8'b01011000;
		sin[304] <= 8'b01011011;
		sin[305] <= 8'b01011101;
		sin[306] <= 8'b01011111;
		sin[307] <= 8'b01100010;
		sin[308] <= 8'b01100100;
		sin[309] <= 8'b01100111;
		sin[310] <= 8'b01101001;
		sin[311] <= 8'b01101100;
		sin[312] <= 8'b01101110;
		sin[313] <= 8'b01110001;
		sin[314] <= 8'b01110011;
		sin[315] <= 8'b01110110;
		sin[316] <= 8'b01111000;
		sin[317] <= 8'b01111011;
		sin[318] <= 8'b01111101;
	 end
	 
    //=======================================================
    //  Structural coding
    //=======================================================
	 always @(posedge clk) begin
		q <= sin[addr];
	 end
	 
endmodule